library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity writer is
port (	
		regnum : IN STD_LOGIC_VECTOR(4 downto 0)
		

);
end writer;

architecture Behavioral of writer is
begin

end architecture;